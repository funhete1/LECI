library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity CmpN is
	generic(N : natural := 8);
	port( input0 : in std_logic_vector(N-1 downto 0);
			input1 : in std_logic_vector(N-1 downto 0);
			equal  : out std_logic;
			notEqual: out std_logic;
			ltSigned : out std_logic;
			ltUnsigned : out std_logic);
end CmpN;


architecture Behavioral of CmpN is 
begin 
	equal <= '1' when (input0 = input1) else '0';
	
	notEqual <= '1' when (input0 /= input1) else '0';
	
	ltSigned <= '1' when (signed(input0) < signed(input1)) else '0';
 
	ltUnsigned <= '1' when (unsigned(input0) < unsigned(input1)) else '0';
end Behavioral; 
						